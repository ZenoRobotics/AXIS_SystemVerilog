
`ifndef _rx_tx_axis_parameters_vh_
`define _rx_tx_axis_parameters_vh_
// Indexes for the lane #'s based on their purpose
parameter LANE_CONTROLLER = 0;
parameter LANE_OUTBOUND = 1;

// Global Variables
parameter NUM_RX_LANES = 2;
parameter NUM_TX_LANES = 2;

`endif